library verilog;
use verilog.vl_types.all;
entity d1s4392 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : out    vl_logic
    );
end d1s4392;
