library verilog;
use verilog.vl_types.all;
entity d1s4812tb is
end d1s4812tb;
